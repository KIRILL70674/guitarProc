module marsohodAudioFPGA();

endmodule:marsohodAudioFPGA