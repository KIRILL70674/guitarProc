module marsohodAudioFPGA();
// test comment
endmodule:marsohodAudioFPGA